// =====================================================================
// Module Name : Initial Permutation Table
// Date : 19/10/2024
// Description : Cryptographic Accelerator
// =====================================================================

module initial_perm(
    input [63:0] data_in,
    output [63:0] out
);
    function [63:0]	IEX;
		input [63:0] D;
		begin	
			IEX[63] = D[64-58];
			IEX[62] = D[64-50];
			IEX[61] = D[64-42];
			IEX[60] = D[64-34];
			IEX[59] = D[64-26];
			IEX[58] = D[64-18];
			IEX[57] = D[64-10];
			IEX[56] = D[64- 2];		
			IEX[55] = D[64-60];
			IEX[54] = D[64-52];
			IEX[53] = D[64-44];
			IEX[52] = D[64-36];
			IEX[51] = D[64-28];
			IEX[50] = D[64-20];
			IEX[49] = D[64-12];
			IEX[48] = D[64- 4];
			IEX[47] = D[64-62];
			IEX[46] = D[64-54];
			IEX[45] = D[64-46];
			IEX[44] = D[64-38];
			IEX[43] = D[64-30];
			IEX[42] = D[64-22];
			IEX[41] = D[64-14];
			IEX[40] = D[64- 6];
			IEX[39] = D[64-64];
			IEX[38] = D[64-56];
			IEX[37] = D[64-48];
			IEX[36] = D[64-40];
			IEX[35] = D[64-32];
			IEX[34] = D[64-24];
			IEX[33] = D[64-16];
			IEX[32] = D[64- 8];
			IEX[31] = D[64-57];
			IEX[30] = D[64-49];
			IEX[29] = D[64-41];
			IEX[28] = D[64-33];
			IEX[27] = D[64-25];
			IEX[26] = D[64-17];
			IEX[25] = D[64- 9];
			IEX[24] = D[64- 1];
			IEX[23] = D[64-59];
			IEX[22] = D[64-51];
			IEX[21] = D[64-43];
			IEX[20] = D[64-35];
			IEX[19] = D[64-27];
			IEX[18] = D[64-19];
			IEX[17] = D[64-11];
			IEX[16] = D[64- 3];
			IEX[15] = D[64-61];
			IEX[14] = D[64-53];
			IEX[13] = D[64-45];
			IEX[12] = D[64-37];
			IEX[11] = D[64-29];
			IEX[10] = D[64-21];
			IEX[ 9] = D[64-13];
			IEX[ 8] = D[64- 5];		
			IEX[ 7] = D[64-63];
			IEX[ 6] = D[64-55];
			IEX[ 5] = D[64-47];
			IEX[ 4] = D[64-39];
			IEX[ 3] = D[64-31];
			IEX[ 2] = D[64-23];
			IEX[ 1] = D[64-15];
			IEX[ 0] = D[64- 7];					
		end
	endfunction

    assign out = IEX(data_in);
    
endmodule