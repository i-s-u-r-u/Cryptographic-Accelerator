// =====================================================================
// Module Name : Final Permutation Table
// Date : 19/10/2024
// Description : Cryptographic Accelerator
// =====================================================================

module final_perm(
    input [63:0] data_in,
    output [63:0] out
);
    function [63:0]	LEX;
		input [63:0] D;
		begin	
			LEX[63] = D[64-40];
			LEX[62] = D[64- 8];
			LEX[61] = D[64-48];
			LEX[60] = D[64-16];
			LEX[59] = D[64-56];
			LEX[58] = D[64-24];
			LEX[57] = D[64-64];
			LEX[56] = D[64-32];		
			LEX[55] = D[64-39];
			LEX[54] = D[64- 7];
			LEX[53] = D[64-47];
			LEX[52] = D[64-15];
			LEX[51] = D[64-55];
			LEX[50] = D[64-23];
			LEX[49] = D[64-63];
			LEX[48] = D[64-31];
			LEX[47] = D[64-38];
			LEX[46] = D[64- 6];
			LEX[45] = D[64-46];
			LEX[44] = D[64-14];
			LEX[43] = D[64-54];
			LEX[42] = D[64-22];
			LEX[41] = D[64-62];
			LEX[40] = D[64-30];
			LEX[39] = D[64-37];
			LEX[38] = D[64- 5];
			LEX[37] = D[64-45];
			LEX[36] = D[64-13];
			LEX[35] = D[64-53];
			LEX[34] = D[64-21];
			LEX[33] = D[64-61];
			LEX[32] = D[64-29];
			LEX[31] = D[64-36];
			LEX[30] = D[64- 4];
			LEX[29] = D[64-44];
			LEX[28] = D[64-12];
			LEX[27] = D[64-52];
			LEX[26] = D[64-20];
			LEX[25] = D[64-60];
			LEX[24] = D[64-28];
			LEX[23] = D[64-35];
			LEX[22] = D[64- 3];
			LEX[21] = D[64-43];
			LEX[20] = D[64-11];
			LEX[19] = D[64-51];
			LEX[18] = D[64-19];
			LEX[17] = D[64-59];
			LEX[16] = D[64-27];
			LEX[15] = D[64-34];
			LEX[14] = D[64- 2];
			LEX[13] = D[64-42];
			LEX[12] = D[64-10];
			LEX[11] = D[64-50];
			LEX[10] = D[64-18];
			LEX[ 9] = D[64-58];
			LEX[ 8] = D[64-26];		
			LEX[ 7] = D[64-33];
			LEX[ 6] = D[64- 1];
			LEX[ 5] = D[64-41];
			LEX[ 4] = D[64- 9];
			LEX[ 3] = D[64-49];
			LEX[ 2] = D[64-17];
			LEX[ 1] = D[64-57];
			LEX[ 0] = D[64-25];					
		end
	endfunction

    assign out = LEX(data_in);
    
endmodule